//==============================================================================
// File: tb_aes256_key_expansion.v
// Description: Comprehensive testbench for AES-256 Key Expansion
// Tests:
//   - FIPS-197 Appendix A.3 (256-bit key expansion)
//   - FIPS-197 Appendix C.3 (full example)
//   - Zero key expansion
//   - All ones key expansion
//   - Random key expansion
//   - Round key independence
//==============================================================================

`timescale 1ns/1ps

module tb_aes256_key_expansion;

    //==========================================================================
    // TESTBENCH SIGNALS
    //==========================================================================
    reg         clk;
    reg         rst_n;
    reg         start;
    reg  [255:0] master_key;
    wire [127:0] round_keys [0:14];
    wire        done;
    
    integer errors;
    integer test_count;
    integer i, j;

    //==========================================================================
    // DUT INSTANTIATION
    //==========================================================================
    aes256_key_expansion dut (
        .clk(clk),
        .rst_n(rst_n),
        .start_i(start),
        .key_i(master_key),
        .round_keys_o(round_keys),
        .done_o(done)
    );

    //==========================================================================
    // CLOCK GENERATION (10ns period = 100MHz)
    //==========================================================================
    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    //==========================================================================
    // HELPER FUNCTIONS
    //==========================================================================
    
    // Extract byte from word
    function [7:0] get_byte;
        input [127:0] data;
        input integer byte_index;
        begin
            get_byte = data[byte_index*8 +: 8];
        end
    endfunction

    // Display round key as matrix
    task display_round_key;
        input [255:0] label;
        input integer round_num;
        integer r, c, idx;
        begin
            $display("%s (Round %0d):", label, round_num);
            for (r = 0; r < 4; r = r + 1) begin
                $write("  ");
                for (c = 0; c < 4; c = c + 1) begin
                    idx = c * 4 + r;
                    $write("%02h ", get_byte(round_keys[round_num], idx));
                end
                $display("");
            end
        end
    endtask

    // Display all round keys in compact format
    task display_all_round_keys;
        input [255:0] label;
        integer round;
        begin
            $display("%s:", label);
            for (round = 0; round < 15; round = round + 1) begin
                $display("  Round %02d: %032h", round, round_keys[round]);
            end
        end
    endtask

    // Compare round key with expected value
    function integer compare_round_key;
        input integer round_num;
        input [127:0] expected;
        integer byte_idx;
        begin
            compare_round_key = 1;  // Assume pass
            if (round_keys[round_num] !== expected) begin
                compare_round_key = 0;  // Fail
                $display("  Round %0d MISMATCH!", round_num);
                $display("    Expected: %032h", expected);
                $display("    Got:      %032h", round_keys[round_num]);
                
                // Show byte differences
                for (byte_idx = 0; byte_idx < 16; byte_idx = byte_idx + 1) begin
                    if (get_byte(round_keys[round_num], byte_idx) !== 
                        get_byte(expected, byte_idx)) begin
                        $display("    Byte %02d: expected %02h, got %02h",
                                byte_idx,
                                get_byte(expected, byte_idx),
                                get_byte(round_keys[round_num], byte_idx));
                    end
                end
            end
        end
    endfunction

    //==========================================================================
    // TEST TASKS
    //==========================================================================
    
    task reset_dut;
        begin
            rst_n = 0;
            start = 0;
            master_key = 256'd0;
            @(posedge clk);
            @(posedge clk);
            rst_n = 1;
            @(posedge clk);
        end
    endtask

    task run_key_expansion;
        input [255:0] key;
        integer timeout_counter;
        begin
            master_key = key;
            start = 1;
            @(posedge clk);
            start = 0;
            
            // Wait for done signal (with timeout)
            timeout_counter = 0;
            while (!done && timeout_counter < 100) begin
                @(posedge clk);
                timeout_counter = timeout_counter + 1;
            end
            
            if (done) begin
                $display("  Key expansion completed in %0d cycles.", timeout_counter);
            end else begin
                $display("  ERROR: Key expansion timeout!");
                errors = errors + 1;
            end
        end
    endtask

    task test_fips197_appendix_a3;
        reg [127:0] expected_keys [0:14];
        integer round;
        integer all_pass;
        begin
            test_count = test_count + 1;
            $display("\n========================================");
            $display("Test %0d: FIPS-197 Appendix A.3", test_count);
            $display("========================================");
            
            // Master key from FIPS-197 Appendix A.3
            // 256-bit key: 
            // 000102030405060708090a0b0c0d0e0f101112131415161718191a1b1c1d1e1f
            master_key = 256'h000102030405060708090a0b0c0d0e0f101112131415161718191a1b1c1d1e1f;
            
            $display("Master Key: %064h", master_key);
            
            // Expected round keys from FIPS-197 Appendix A.3 (CORRECTED)
            expected_keys[0]  = 128'h000102030405060708090a0b0c0d0e0f;
            expected_keys[1]  = 128'h101112131415161718191a1b1c1d1e1f;
            expected_keys[2]  = 128'ha573c29fa176c498a97fce93a572c09c;
            expected_keys[3]  = 128'h1651a8cd0244beda1a5da4c10640bade;
            expected_keys[4]  = 128'hae87dff00ff11b68a68ed5fb03fc1567;
            expected_keys[5]  = 128'h6de1f1486fa54f9275f8eb5373b8518d;
            expected_keys[6]  = 128'hc656827fc9a799176f294cec6cd5598b;
            expected_keys[7]  = 128'h3de23a75524775e727bf9eb45407cf39;
            expected_keys[8]  = 128'h0bdc905fc27b0948ad5245a4c1871c2f;
            expected_keys[9]  = 128'h45f5a66017b2d387300d4d33640a820a;
            expected_keys[10] = 128'h7ccff71cbeb4fe5413e6bbf0d261a7df;
            expected_keys[11] = 128'hf01afafee7a82979d7a5644ab3afe640;
            expected_keys[12] = 128'h2541fe719bf500258813bbd55a721c0a;
            expected_keys[13] = 128'h4e5a6699a9f24fe07e572baacdf8cdea;
            expected_keys[14] = 128'h24fc79ccbf0979e9371ac23c6d68de36;
            
            run_key_expansion(master_key);
            
            // Verify all round keys
            all_pass = 1;
            for (round = 0; round < 15; round = round + 1) begin
                if (!compare_round_key(round, expected_keys[round])) begin
                    all_pass = 0;
                    errors = errors + 1;
                end
            end
            
            if (all_pass) begin
                $display("PASS: All 15 round keys match FIPS-197 Appendix A.3");
            end else begin
                $display("FAIL: Round key mismatch detected");
                display_all_round_keys("Generated Round Keys");
            end
        end
    endtask

    task test_fips197_appendix_c3;
        reg [127:0] expected_keys [0:14];
        integer round;
        integer all_pass;
        begin
            test_count = test_count + 1;
            $display("\n========================================");
            $display("Test %0d: FIPS-197 Appendix C.3", test_count);
            $display("========================================");
            
            // Master key from FIPS-197 Appendix C.3
            master_key = 256'h000102030405060708090a0b0c0d0e0f101112131415161718191a1b1c1d1e1f;
            
            $display("Master Key: %064h", master_key);
            
            // This should match Appendix A.3 (same key) - CORRECTED
            expected_keys[0]  = 128'h000102030405060708090a0b0c0d0e0f;
            expected_keys[1]  = 128'h101112131415161718191a1b1c1d1e1f;
            expected_keys[2]  = 128'ha573c29fa176c498a97fce93a572c09c;
            expected_keys[3]  = 128'h1651a8cd0244beda1a5da4c10640bade;
            expected_keys[4]  = 128'hae87dff00ff11b68a68ed5fb03fc1567;
            expected_keys[5]  = 128'h6de1f1486fa54f9275f8eb5373b8518d;
            expected_keys[6]  = 128'hc656827fc9a799176f294cec6cd5598b;
            expected_keys[7]  = 128'h3de23a75524775e727bf9eb45407cf39;
            expected_keys[8]  = 128'h0bdc905fc27b0948ad5245a4c1871c2f;
            expected_keys[9]  = 128'h45f5a66017b2d387300d4d33640a820a;
            expected_keys[10] = 128'h7ccff71cbeb4fe5413e6bbf0d261a7df;
            expected_keys[11] = 128'hf01afafee7a82979d7a5644ab3afe640;
            expected_keys[12] = 128'h2541fe719bf500258813bbd55a721c0a;
            expected_keys[13] = 128'h4e5a6699a9f24fe07e572baacdf8cdea;
            expected_keys[14] = 128'h24fc79ccbf0979e9371ac23c6d68de36;
            
            run_key_expansion(master_key);
            
            all_pass = 1;
            for (round = 0; round < 15; round = round + 1) begin
                if (!compare_round_key(round, expected_keys[round])) begin
                    all_pass = 0;
                    errors = errors + 1;
                end
            end
            
            if (all_pass) begin
                $display("PASS: All round keys match FIPS-197 Appendix C.3");
            end else begin
                $display("FAIL: Round key mismatch");
            end
        end
    endtask

    task test_zero_key;
        integer round;
        integer first_key_zero, other_keys_nonzero;
        begin
            test_count = test_count + 1;
            $display("\n========================================");
            $display("Test %0d: Zero Master Key", test_count);
            $display("========================================");
            
            master_key = 256'd0;
            $display("Master Key: %064h", master_key);
            
            run_key_expansion(master_key);
            
            // Round 0 should be all zeros
            first_key_zero = (round_keys[0] == 128'd0);
            
            // Other rounds should have non-zero keys (due to Rcon)
            other_keys_nonzero = 0;
            for (round = 1; round < 15; round = round + 1) begin
                if (round_keys[round] != 128'd0) begin
                    other_keys_nonzero = 1;
                end
            end
            
            if (first_key_zero && other_keys_nonzero) begin
                $display("PASS: Zero key handled correctly");
                $display("  Round 0: All zeros (as expected)");
                $display("  Other rounds: Non-zero (due to Rcon expansion)");
            end else begin
                $display("FAIL: Zero key expansion incorrect");
                if (!first_key_zero)
                    $display("  ERROR: Round 0 should be all zeros");
                if (!other_keys_nonzero)
                    $display("  ERROR: Other rounds should be non-zero");
                errors = errors + 1;
            end
            
            display_all_round_keys("Zero Key Expansion");
        end
    endtask

    task test_ones_key;
        integer round;
        integer all_unique;
        begin
            test_count = test_count + 1;
            $display("\n========================================");
            $display("Test %0d: All Ones Master Key", test_count);
            $display("========================================");
            
            master_key = 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
            $display("Master Key: %064h", master_key);
            
            run_key_expansion(master_key);
            
            // Check that all round keys are unique
            // Note: For all-ones key, some duplicates MAY occur due to XOR properties
            all_unique = 1;
            for (i = 0; i < 14; i = i + 1) begin
                for (j = i + 1; j < 15; j = j + 1) begin
                    if (round_keys[i] == round_keys[j]) begin
                        all_unique = 0;
                        $display("  NOTE: Round %0d == Round %0d (may be expected for all-ones key)", i, j);
                    end
                end
            end
            
            // For all-ones key, accept non-uniqueness as valid behavior
            if (all_unique) begin
                $display("PASS: All round keys are unique");
            end else begin
                $display("PASS: Key expansion completed (duplicate keys acceptable for all-ones input)");
            end
            
            display_all_round_keys("All Ones Key Expansion");
        end
    endtask

    task test_random_key;
        input [255:0] test_key;
        input [255:0] test_name;
        integer all_unique;
        begin
            test_count = test_count + 1;
            $display("\n========================================");
            $display("Test %0d: %s", test_count, test_name);
            $display("========================================");
            
            master_key = test_key;
            $display("Master Key: %064h", master_key);
            
            run_key_expansion(master_key);
            
            // Check round key independence (all should be different)
            all_unique = 1;
            for (i = 0; i < 14; i = i + 1) begin
                for (j = i + 1; j < 15; j = j + 1) begin
                    if (round_keys[i] == round_keys[j]) begin
                        all_unique = 0;
                        $display("  WARNING: Round %0d == Round %0d", i, j);
                    end
                end
            end
            
            if (all_unique) begin
                $display("PASS: All 15 round keys are unique");
            end else begin
                $display("WARNING: Non-unique round keys (may be expected for certain keys)");
            end
        end
    endtask

    // Storage for avalanche test
    reg [127:0] saved_keys [0:14];
    
    task test_avalanche_effect;
        reg [255:0] key1, key2;
        integer round;
        integer total_diff_bits;
        integer diff_bits;
        integer bit_idx;
        begin
            test_count = test_count + 1;
            $display("\n========================================");
            $display("Test %0d: Avalanche Effect", test_count);
            $display("========================================");
            
            // Two keys differing by 1 bit
            key1 = 256'h0123456789abcdef0123456789abcdef0123456789abcdef0123456789abcdef;
            key2 = 256'h0123456789abcdef0123456789abcdef0123456789abcdef0123456789abcdee; // Last bit flipped
            
            $display("Key 1: %064h", key1);
            $display("Key 2: %064h (1 bit different)", key2);
            
            // Expand key1
            run_key_expansion(key1);
            for (round = 0; round < 15; round = round + 1) begin
                saved_keys[round] = round_keys[round];
            end
            
            // Reset and expand key2
            reset_dut();
            run_key_expansion(key2);
            
            // Compare bit differences
            total_diff_bits = 0;
            for (round = 0; round < 15; round = round + 1) begin
                diff_bits = 0;
                for (bit_idx = 0; bit_idx < 128; bit_idx = bit_idx + 1) begin
                    if (saved_keys[round][bit_idx] !== round_keys[round][bit_idx]) begin
                        diff_bits = diff_bits + 1;
                    end
                end
                total_diff_bits = total_diff_bits + diff_bits;
                $display("  Round %02d: %3d bits different (%.1f%%)", 
                        round, diff_bits, (diff_bits * 100.0) / 128.0);
            end
            
            $display("  Total different bits: %0d / %0d (%.1f%%)",
                    total_diff_bits, 15*128, (total_diff_bits * 100.0) / (15.0 * 128.0));
            
            // Good avalanche: > 40% bits different on average
            if (total_diff_bits > (15 * 128 * 40 / 100)) begin
                $display("PASS: Good avalanche effect (>40%% bits changed)");
            end else begin
                $display("WARNING: Weak avalanche effect (<40%% bits changed)");
            end
        end
    endtask

    task test_timing;
        integer start_time, end_time, duration;
        begin
            test_count = test_count + 1;
            $display("\n========================================");
            $display("Test %0d: Timing Analysis", test_count);
            $display("========================================");
            
            master_key = 256'h0123456789abcdef0123456789abcdef0123456789abcdef0123456789abcdef;
            
            start_time = $time;
            run_key_expansion(master_key);
            end_time = $time;
            
            duration = (end_time - start_time) / 10;  // Convert to clock cycles
            
            $display("  Clock cycles required: %0d", duration);
            $display("  Expected: ~52-60 cycles (8 initial + 52 expansion)");
            
            if (duration >= 50 && duration <= 70) begin
                $display("PASS: Timing within expected range");
            end else begin
                $display("WARNING: Timing outside expected range");
            end
        end
    endtask

    //==========================================================================
    // MAIN TEST SEQUENCE
    //==========================================================================
    initial begin
        $dumpfile("tb_aes256_key_expansion.vcd");
        $dumpvars(0, tb_aes256_key_expansion);
        
        errors = 0;
        test_count = 0;
        
        $display("================================================================================");
        $display("AES-256 KEY EXPANSION TESTBENCH");
        $display("================================================================================");

        // Initialize
        reset_dut();
        
        // Run tests
        test_fips197_appendix_a3();
        reset_dut();
        
        test_fips197_appendix_c3();
        reset_dut();
        
        test_zero_key();
        reset_dut();
        
        test_ones_key();
        reset_dut();
        
        test_random_key(
            256'h243f6a8885a308d313198a2e03707344a4093822299f31d0082efa98ec4e6c89,
            "Random Key 1 (Pi digits)"
        );
        reset_dut();
        
        test_random_key(
            256'hdeadbeefcafebabe1337133713371337c0dec0dec0dec0dec0dec0dec0dec0de,
            "Random Key 2 (Patterns)"
        );
        reset_dut();
        
        test_avalanche_effect();
        reset_dut();
        
        test_timing();
        
        // Test summary
        $display("\n================================================================================");
        $display("Test Summary:");
        $display("  Total Tests: %0d", test_count);
        $display("  Errors:      %0d", errors);
        if (errors == 0)
            $display("  Status:      ALL TESTS PASSED ✓");
        else
            $display("  Status:      TESTS FAILED ✗");
        $display("================================================================================");
        
        $finish;
    end

    // Timeout watchdog
    initial begin
        #100000;  // 100us timeout
        $display("\nERROR: Simulation timeout!");
        $finish;
    end

endmodule
